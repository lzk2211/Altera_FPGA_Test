library verilog;
use verilog.vl_types.all;
entity u_addr_vlg_vec_tst is
end u_addr_vlg_vec_tst;
