library verilog;
use verilog.vl_types.all;
entity u_addr_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end u_addr_vlg_sample_tst;
