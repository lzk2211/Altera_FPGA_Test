library verilog;
use verilog.vl_types.all;
entity aa_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end aa_vlg_sample_tst;
