library verilog;
use verilog.vl_types.all;
entity smg_display_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end smg_display_vlg_sample_tst;
