library verilog;
use verilog.vl_types.all;
entity switch_scoure_vlg_check_tst is
    port(
        outp            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end switch_scoure_vlg_check_tst;
