library verilog;
use verilog.vl_types.all;
entity bjq_vlg_vec_tst is
end bjq_vlg_vec_tst;
