library verilog;
use verilog.vl_types.all;
entity tst2_vlg_vec_tst is
end tst2_vlg_vec_tst;
