library verilog;
use verilog.vl_types.all;
entity smg_display1_vlg_vec_tst is
end smg_display1_vlg_vec_tst;
