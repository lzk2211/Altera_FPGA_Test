library verilog;
use verilog.vl_types.all;
entity tst1_38_vlg_vec_tst is
end tst1_38_vlg_vec_tst;
