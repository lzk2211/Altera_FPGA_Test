library verilog;
use verilog.vl_types.all;
entity tst1_38 is
    port(
        Y1              : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        Y2              : out    vl_logic;
        Y4              : out    vl_logic;
        Y3              : out    vl_logic;
        Y5              : out    vl_logic;
        Y6              : out    vl_logic;
        Y7              : out    vl_logic;
        Y0              : out    vl_logic
    );
end tst1_38;
