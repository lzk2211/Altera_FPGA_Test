library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity cnt_time is
port(nreset: in std_logic;
	  clk: in std_logic;
	  
	  count_sec: out std_logic_vector(3 downto 0);
	  LED8s: out std_logic_vector(7 downto 0);
	  SEL: out std_logic_vector(2 downto 0)
	  );
end;

architecture behav of cnt_time is
signal count: std_logic_vector(3 downto 0) := "0000";
signal SE: std_logic_vector(2 downto 0) := "000";
begin
	process(nreset, clk)
	begin
		if nreset = '0' then
			count <= "0000";
			SE <= "111";
			
		elsif clk' event and clk = '1' then
			if count >= "1001" then
				count <= "0000";
			else
				count <= count + 1;
			end if;
			
			SE <= SE + 1;
			
		end if;
	end process;
	
	count_sec <= count;
	
	LED8s <= "00111111" when count = "0000" else
				"00000110" when count = "0001" else
				"01011011" when count = "0010" else
				"01001111" when count = "0011" else
				"01100110" when count = "0100" else
				"01101101" when count = "0101" else
				"01111101" when count = "0110" else
				"00000111" when count = "0111" else
				"01111111" when count = "1000" else
				"01101111" when count = "1001" else
				"00000000";
				
	SEL <= SE;	
end;