library verilog;
use verilog.vl_types.all;
entity switch_scoure_vlg_vec_tst is
end switch_scoure_vlg_vec_tst;
