library verilog;
use verilog.vl_types.all;
entity count_add_vlg_vec_tst is
end count_add_vlg_vec_tst;
