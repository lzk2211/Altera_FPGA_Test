library verilog;
use verilog.vl_types.all;
entity aa_vlg_vec_tst is
end aa_vlg_vec_tst;
